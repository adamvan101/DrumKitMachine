kick-tape
kick-tape
snare-808
snare-808
hihat-808
hihat-808
tom-acoustic02
clap-808
tom-acoustic01
clap-808
tom-808
tom-acoustic01
crash-tape
tom-acoustic02
ride-acoustic01
clap-808
crash-acoustic
clap-808
